package waveform_lut_pkg is
type t_sine_array is array (0 to 255) of natural;
constant sine_lut : t_sine_array :=
	(8388608,
	8594474,
	8800217,
	9005712,
	9210835,
	9415463,
	9619472,
	9822740,
	10025144,
	10226562,
	10426873,
	10625956,
	10823692,
	11019961,
	11214644,
	11407626,
	11598789,
	11788018,
	11975199,
	12160220,
	12342970,
	12523337,
	12701214,
	12876493,
	13049068,
	13218836,
	13385695,
	13549544,
	13710284,
	13867818,
	14022052,
	14172892,
	14320249,
	14464032,
	14604156,
	14740535,
	14873089,
	15001736,
	15126400,
	15247006,
	15363480,
	15475752,
	15583756,
	15687426,
	15786699,
	15881516,
	15971819,
	16057554,
	16138670,
	16215118,
	16286851,
	16353827,
	16416004,
	16473347,
	16525819,
	16573390,
	16616030,
	16653715,
	16686421,
	16714129,
	16736822,
	16754486,
	16767111,
	16774689,
	16777215,
	16774689,
	16767111,
	16754486,
	16736822,
	16714129,
	16686421,
	16653715,
	16616030,
	16573390,
	16525819,
	16473347,
	16416004,
	16353827,
	16286851,
	16215118,
	16138670,
	16057554,
	15971819,
	15881516,
	15786699,
	15687426,
	15583756,
	15475752,
	15363480,
	15247006,
	15126400,
	15001736,
	14873089,
	14740535,
	14604156,
	14464032,
	14320249,
	14172892,
	14022052,
	13867818,
	13710284,
	13549544,
	13385695,
	13218836,
	13049068,
	12876493,
	12701214,
	12523337,
	12342970,
	12160220,
	11975199,
	11788018,
	11598789,
	11407626,
	11214644,
	11019961,
	10823692,
	10625956,
	10426873,
	10226562,
	10025144,
	9822740,
	9619472,
	9415463,
	9210835,
	9005712,
	8800217,
	8594474,
	8388608,
	8182741,
	7976998,
	7771503,
	7566380,
	7361752,
	7157743,
	6954475,
	6752071,
	6550653,
	6350342,
	6151259,
	5953523,
	5757254,
	5562571,
	5369589,
	5178426,
	4989197,
	4802016,
	4616995,
	4434245,
	4253878,
	4076001,
	3900722,
	3728147,
	3558379,
	3391520,
	3227671,
	3066931,
	2909397,
	2755163,
	2604323,
	2456966,
	2313183,
	2173059,
	2036680,
	1904126,
	1775479,
	1650815,
	1530209,
	1413735,
	1301463,
	1193459,
	1089789,
	990516,
	895699,
	805396,
	719661,
	638545,
	562097,
	490364,
	423388,
	361211,
	303868,
	251396,
	203825,
	161185,
	123500,
	90794,
	63086,
	40393,
	22729,
	10104,
	2526,
	0,
	2526,
	10104,
	22729,
	40393,
	63086,
	90794,
	123500,
	161185,
	203825,
	251396,
	303868,
	361211,
	423388,
	490364,
	562097,
	638545,
	719661,
	805396,
	895699,
	990516,
	1089789,
	1193459,
	1301463,
	1413735,
	1530209,
	1650815,
	1775479,
	1904126,
	2036680,
	2173059,
	2313183,
	2456966,
	2604323,
	2755163,
	2909397,
	3066931,
	3227671,
	3391520,
	3558379,
	3728147,
	3900722,
	4076001,
	4253878,
	4434245,
	4616995,
	4802016,
	4989197,
	5178426,
	5369589,
	5562571,
	5757254,
	5953523,
	6151259,
	6350342,
	6550653,
	6752071,
	6954475,
	7157743,
	7361752,
	7566380,
	7771503,
	7976998,
	8182741);

end package waveform_lut_pkg;

package body waveform_lut_pkg is

end package body waveform_lut_pkg;
